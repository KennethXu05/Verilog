module alu74181_alu74182_16bit_tb();
    reg [15:0] A;
    reg [15:0] B;
    reg Cin;
    wire [15:0] S;

    cla_16bit u_cla_16bit(
        .A  (A),
        .B  (B),
        .Cin(Cin),
        .S  (S)
    );

    initial begin
        A = 16'b0000_0000_0000_0000; B = 16'b0000_0000_0000_0000; Cin = 1'b0;
        #10 A = 16'b0000_0000_0000_0001; B = 16'b0000_0000_0000_0010; Cin = 1'b0;
        #10 A = 16'b0000_0000_0000_0011; B = 16'b0000_0000_0000_0100; Cin = 1'b0;
        #10 A = 16'b0000_0000_0000_0101; B = 16'b0000_0000_0000_0110; Cin = 1'b0;
        #10 A = 16'b0000_0000_0000_0111; B = 16'b0000_0000_0000_1000; Cin = 1'b0;
        #10 A = 16'b0000_0000_0000_1001; B = 16'b0000_0000_0000_1010; Cin = 1'b0;
        #10 A = 16'b0000_0000_0000_1011; B = 16'b0000_0000_0000_1100; Cin = 1'b0;
        #10 A = 16'b0000_0000_0000_1101; B = 16'b0000_0000_0000_1110; Cin = 1'b0;
        #10 A = 16'b0000_0000_0000_1111; B = 16'b0000_0000_0000_0001; Cin = 1'b0;
        #10 A = 16'b1111_1111_1111_1111; B = 16'b1111_1111_1111_1111; Cin = 1'b1;
        #10 $stop;
    end
endmodule